LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
-----------------------------------------------------
ENTITY DPLDRV IS
	PORT (   CLK50M		:	IN		STD_LOGIC;
				DIGITO0		:	IN		INTEGER RANGE 0 TO 15;
				DIGITO1		:	IN		INTEGER RANGE 0 TO 15;
				DIGITO2		:	IN		INTEGER RANGE 0 TO 15;
				DIGITO3		:	IN		INTEGER RANGE 0 TO 15;
				DPL_ENABLE	:	OUT 	STD_LOGIC_VECTOR (3  DOWNTO 0);
				DPL_SEG		:	OUT 	STD_LOGIC_VECTOR	(6  DOWNTO 0)
-----------------------------------------------------------------
         );
END DPLDRV;
--------------------------
ARCHITECTURE BEHAVIORAL OF DPLDRV IS
SIGNAL	DIGITO		:	INTEGER RANGE 0 TO 15:=0;
SIGNAL	POS_DISPLAY	:	INTEGER RANGE 0 TO 3:=0;
SIGNAL	DELAY			:	STD_LOGIC_VECTOR (13  DOWNTO 0);
BEGIN
	DPL_ENABLE	<=	"1110"	WHEN	(POS_DISPLAY = 0)	ELSE
						"1101"	WHEN	(POS_DISPLAY = 1)	ELSE
						"1011"	WHEN	(POS_DISPLAY = 2)	ELSE
						"0111";
	DIGITO		<=	DIGITO0	WHEN	(POS_DISPLAY = 0)	ELSE
						DIGITO1	WHEN	(POS_DISPLAY = 1)	ELSE
						DIGITO2	WHEN	(POS_DISPLAY = 2)	ELSE
						DIGITO3;
	DPL_SEG		<=	"0000001"	WHEN	(DIGITO=0)	ELSE
						"1001111"	WHEN	(DIGITO=1)	ELSE
						"0010010"	WHEN	(DIGITO=2)	ELSE
						"0000110"	WHEN	(DIGITO=3)	ELSE
						"1001100"	WHEN	(DIGITO=4)	ELSE
						"0100100"	WHEN	(DIGITO=5)	ELSE
						"0100000"	WHEN	(DIGITO=6)	ELSE
						"0001111"	WHEN	(DIGITO=7)	ELSE
						"0000000"	WHEN	(DIGITO=8)	ELSE
						"0000100"	WHEN	(DIGITO=9)	ELSE
						"1111111";
	PROCESS (CLK50M)
	BEGIN
		IF (CLK50M'EVENT AND CLK50M='1') THEN
			DELAY	<=	DELAY+1;
			IF ( DELAY="11111111111111" ) THEN
				POS_DISPLAY	<=	POS_DISPLAY+1;
			END IF;
		END IF;
	END PROCESS;
END BEHAVIORAL;