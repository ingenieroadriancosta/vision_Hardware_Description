LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
-----------------------------------------------------
ENTITY BYTE2BCD IS
	PORT (   BYTE2IN 		:	IN    NATURAL RANGE 0 TO 31;
				DIGITO0   	:	OUT   NATURAL RANGE 0 TO 15;
				DIGITO1   	:	OUT   NATURAL RANGE 0 TO 15
-----------------------------------------------------------------
         );
END BYTE2BCD;
-----------------------------------------------------
ARCHITECTURE BEHAVIORAL OF BYTE2BCD IS

SIGNAL	DU1			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU2			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU3			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );



SIGNAL	DD0			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );



SIGNAL	BYTE			:	STD_LOGIC_VECTOR( 4 DOWNTO 0 );


BEGIN
	BYTE	<=	CONV_STD_LOGIC_VECTOR( BYTE2IN , 5 );
	--UNIDADES.

	DU1	<=	'0'&BYTE(4 DOWNTO 2)				WHEN	( ('0'&BYTE(4 DOWNTO 2))<5 )	ELSE
				'0'&BYTE(4 DOWNTO 2)+3;
	DU2	<=	DU1(2 DOWNTO 0)&BYTE(1)	WHEN	( (DU1(2 DOWNTO 0)&BYTE(1))<5 )	ELSE
				DU1(2 DOWNTO 0)&BYTE(1)+3;
	DU3	<=	DU2(2 DOWNTO 0)&BYTE(0);
	
	
	--DECENAS.
	DD0	<=	'0'&'0'&DU1(3)&DU2(3);
	

	DIGITO0	<=	CONV_INTEGER(DU3);
	DIGITO1	<=	CONV_INTEGER(DD0);
--	DIGITO2	<=	CONV_INTEGER(DC0);
--	DIGITO3	<=	CONV_INTEGER(PRBDATA);
END BEHAVIORAL;