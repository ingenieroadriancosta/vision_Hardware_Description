LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE PAQUETE IS


SIGNAL	CLK0DLL		:	STD_LOGIC;
SIGNAL	CLK180DLL	:	STD_LOGIC;
SIGNAL	CLK270DLL	:	STD_LOGIC;
SIGNAL	CLK90DLL	:	STD_LOGIC;
SIGNAL	CLKDVDLL	:	STD_LOGIC;
SIGNAL	LOCKEDDLL	:	STD_LOGIC;




COMPONENT clkDllCtrl IS
  port(ckIn: in std_logic;
       ckOut: inout std_logic
       --ckDivOut: inout std_logic
		 );
END COMPONENT;




COMPONENT USBRECEIVER IS
	PORT(	MCLK			:	IN STD_LOGIC;
			ABORT			:	IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PDB			:	INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			ASTB			:	IN STD_LOGIC;
			DSTB			:	IN STD_LOGIC;
			PWRITE		:	IN STD_LOGIC;
			PWAIT			:	OUT STD_LOGIC;
			
			WORDDATA		:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			PUTDATA		:	OUT BOOLEAN;
			ABORTED		:	OUT BOOLEAN
			);
END COMPONENT;





--SE�ALES PARA LAS ACCIONES DE TECLADO,
SIGNAL	ENABLE_KB	:	BOOLEAN;
SIGNAL	KEY_DOWN		:	BOOLEAN;
SIGNAL	KEY_UP		:	BOOLEAN;
SIGNAL	E0				:	BOOLEAN;
SIGNAL	CTRL			:	BOOLEAN:=FALSE;
SIGNAL	ALT			:	BOOLEAN:=FALSE;
SIGNAL 	RESET			:	BOOLEAN:=FALSE;
SIGNAL 	KBRD_DATA	:	STD_LOGIC_VECTOR (7 DOWNTO 0);

COMPONENT KBRD_PS2 IS
	PORT	(	CLK50M			:	IN  STD_LOGIC;
				KBRD_DATA_PIN 	:	IN  STD_LOGIC;
				KBRD_CLK_PIN	:	IN  STD_LOGIC;
				RESET				:	IN  BOOLEAN;
				KBRD_DATA		:	BUFFER  STD_LOGIC_VECTOR (7 DOWNTO 0);
				ENABLE_KB		:	OUT BOOLEAN;
				KEY_DOWN			:	BUFFER BOOLEAN;
				KEY_UP			:	BUFFER BOOLEAN;
				E0					:	BUFFER BOOLEAN
				
			);
END COMPONENT;





COMPONENT WORD2BCD IS
	PORT (   VARWORD	:	IN    STD_LOGIC_VECTOR (15  DOWNTO 0);
				UNIDAD	:	OUT   STD_LOGIC_VECTOR (3  DOWNTO 0);
				DECENA	:	OUT   STD_LOGIC_VECTOR (3  DOWNTO 0);
				CENTENA	:	OUT   STD_LOGIC_VECTOR (3  DOWNTO 0)
         );
END COMPONENT;



COMPONENT BYTE2BCD IS
	PORT (   BYTE2IN 		:	IN    NATURAL RANGE 0 TO 31;
				DIGITO0   	:	OUT   NATURAL RANGE 0 TO 15;
				DIGITO1   	:	OUT   NATURAL RANGE 0 TO 15
         );
END COMPONENT;




COMPONENT BYTE2BCDALL IS
	PORT (   BYTE    		:	IN    STD_LOGIC_VECTOR (7  DOWNTO 0);
				DIGITO0   	:	OUT   NATURAL RANGE 0 TO 15;
				DIGITO1   	:	OUT   NATURAL RANGE 0 TO 15;
				DIGITO2   	:	OUT   NATURAL RANGE 0 TO 15
-----------------------------------------------------------------
         );
END COMPONENT;



------------------------------------------------------------------------
COMPONENT VGADRVR IS
	PORT( CLK50M		:	IN STD_LOGIC;
			--
			VGA_16_8		:	IN BOOLEAN;
			NORM_NEGA	:	IN BOOLEAN;
			SKD			:	IN BOOLEAN;
			MARK			:	IN BOOLEAN;
			ZOOM			:	IN NATURAL RANGE 0   TO 7;
			COLOR_LETTER:	IN STD_LOGIC_VECTOR (7  DOWNTO 0);
			COLOR_RED	:	IN STD_LOGIC_VECTOR (5  DOWNTO 0);
			COLOR_GREEN	:	IN STD_LOGIC_VECTOR (5  DOWNTO 0);
			COLOR_BLUE	:	IN STD_LOGIC_VECTOR (3  DOWNTO 0);
			--
			MOVE_X		:	IN NATURAL RANGE 0 TO 640:=0;
			MOVE_Y		:	IN NATURAL RANGE 0 TO 480:=0;
			--
			CNT_RAM_POS	:	OUT NATURAL RANGE 0   TO 524287;
			POS_X			:	OUT STD_LOGIC_VECTOR (9  DOWNTO 0);
			POS_Y			:	OUT STD_LOGIC_VECTOR (8  DOWNTO 0);
			--VGA.
			RED			:	OUT STD_LOGIC_VECTOR	(2  DOWNTO 0);
			GRN			:	OUT STD_LOGIC_VECTOR	(2  DOWNTO 0);
			BLUE			:	OUT STD_LOGIC_VECTOR	(1  DOWNTO 0);
			HS				:	OUT STD_LOGIC;
			VS				:	OUT STD_LOGIC
         );
END COMPONENT;












TYPE	MARK	IS	ARRAY	(0 TO 31)	OF	STD_LOGIC_VECTOR (0  TO 127);

CONSTANT	BY_ADRIAN_C_MARK	:	MARK:=(
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11100001111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11000000110001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11000000100011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11001001100100011111111111100111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111",
"10001000000000000111111110000111111100111111111111111111111111111111111111111111111110001001111111111111111111111111111111111111",
"11000011100000001111111100001111111000111111111111111111111111111111111111111111111000111001111111111111111111111111111111111111",
"11000111100000011111110000001111110001111111111100011111111111111111111111111111110001110001111111111111111111100111111111111111",
"11111111111000111111100100011111110011111111111100111111111111111111111111111111100011100011111111111111111111001111111111111111",
"11111111110001111111001100111111100011111111111111111110001111111111111111111111000110000011111111111100111000000111100011111111",
"11111111110011110000011000111100000111000001110001111000001111111100111111111110001100000111100001111100010000001110000011111111",
"11111111110011100000000000010000000110000001100011100000001110000000111111111100011000001110000001111000011100111000000011111111",
"11111111111111000000000000100011001110010011000111000010011100010001111111111100010000011100010001110000011001110000100111111111",
"11111111111111100011100011100100001110100111001111001100011100000001111111111000110001111100110001101100110001100011000111111111",
"11111111111111001111100111100000001001100100001100001000000000000011111111111000111111111000110001000000000000000010000001111111",
"11111111111100011111000001100000000011100001000001000000001100010000111111110000111111100000100001100000110000110000000011100011",
"11111111111100111111000111100010000111100011000011000100011100100001111111110000111111001110001111110001110001110001000111100111",
"11111111111001111111111111111111111111111111111111111111111111111111111111110000111100011111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
);







FUNCTION TO_BIT	(BLIN :	IN BOOLEAN) RETURN STD_LOGIC;
END PAQUETE;



PACKAGE BODY PAQUETE IS

FUNCTION TO_BIT	(BLIN :	IN BOOLEAN) RETURN STD_LOGIC IS
BEGIN
	IF BLIN THEN
		RETURN ('1');
	ELSE
		RETURN ('0');
	END IF;
END TO_BIT;




END PAQUETE;
