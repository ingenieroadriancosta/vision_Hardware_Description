LIBRARY UNISIM;
USE UNISIM.VCOMPONENTS.ALL;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL ;
USE WORK.PAQUETE.ALL;
------------------------------------------------------------------------
ENTITY VGADRVR IS
	PORT( CLK50M		:	IN STD_LOGIC;
			--
			VGA_16_8		:	IN BOOLEAN;
			NORM_NEGA	:	IN BOOLEAN;
			SKD			:	IN BOOLEAN;
			MARK			:	IN	BOOLEAN;
			ZOOM			:	IN NATURAL RANGE 0   TO 7;
			COLOR_LETTER:	IN STD_LOGIC_VECTOR (7  DOWNTO 0);
			COLOR_RED	:	IN STD_LOGIC_VECTOR (5  DOWNTO 0);
			COLOR_GREEN	:	IN STD_LOGIC_VECTOR (5  DOWNTO 0);
			COLOR_BLUE	:	IN STD_LOGIC_VECTOR (3  DOWNTO 0);
			--
			MOVE_X		:	IN NATURAL RANGE 0 TO 640:=0;
			MOVE_Y		:	IN NATURAL RANGE 0 TO 480:=0;
			--
			CNT_RAM_POS	:	OUT NATURAL RANGE 0   TO 524287;
			POS_X			:	OUT STD_LOGIC_VECTOR (9  DOWNTO 0);
			POS_Y			:	OUT STD_LOGIC_VECTOR (8  DOWNTO 0);
			--VGA.
			RED			:	OUT STD_LOGIC_VECTOR	(2  DOWNTO 0);
			GRN			:	OUT STD_LOGIC_VECTOR	(2  DOWNTO 0);
			BLUE			:	OUT STD_LOGIC_VECTOR	(1  DOWNTO 0);
			HS				:	OUT STD_LOGIC;
			VS				:	OUT STD_LOGIC
         );

-- force synthesizer to extract distributed ram for the
-- displayrom signal, and not a block ram, because the block ram
-- is entirely used to store the image.
attribute rom_extract : string;
attribute rom_extract of VGADRVR: entity is "yes";
attribute rom_style : string;
attribute rom_style of VGADRVR: entity is "distributed";

END VGADRVR;

ARCHITECTURE BEHAVIORAL OF VGADRVR IS
SIGNAL	ZERO_COLOR	:	STD_LOGIC_VECTOR (7  DOWNTO 0):="00000000";
SIGNAL	CLK25M		:	STD_LOGIC:='0';
----------------------------------------------------------------------------------------
--SIGNAL	AREA_NEGRA				: BOOLEAN;
--CONTADORES DE BARRIDOS HORIZONTAL Y VERTICAL.
SIGNAL	COUNTER_H		:	STD_LOGIC_VECTOR (9  DOWNTO 0):=(OTHERS=>'0');
SIGNAL	COUNTER_V		:	STD_LOGIC_VECTOR (9  DOWNTO 0):=(OTHERS=>'0');

SIGNAL	COUNTER_H_CUR	:	STD_LOGIC_VECTOR (9  DOWNTO 0);
SIGNAL	COUNTER_V_CUR	:	STD_LOGIC_VECTOR (9  DOWNTO 0);


SIGNAL	POS_X_S			:	STD_LOGIC_VECTOR (9  DOWNTO 0);
SIGNAL	POS_Y_S			:	STD_LOGIC_VECTOR (8  DOWNTO 0);


SIGNAL	COLOR				:	STD_LOGIC_VECTOR (7  DOWNTO 0);
SIGNAL	COLOR_8_BITS	:	STD_LOGIC_VECTOR (7  DOWNTO 0);
SIGNAL	COLOR_16_BITS	:	STD_LOGIC_VECTOR (7  DOWNTO 0);


SIGNAL	VGA_16_8_VECTOR:	STD_LOGIC_VECTOR (7  DOWNTO 0);
--SIGNAL	COMPLETE				:	BOOLEAN:=FALSE;


SIGNAL	TOCOLORRED	:	STD_LOGIC_VECTOR (2  DOWNTO 0);
SIGNAL	TOCOLORGREEN:	STD_LOGIC_VECTOR (2  DOWNTO 0);
SIGNAL	TOCOLORBLUE	:	STD_LOGIC_VECTOR (1  DOWNTO 0);


SIGNAL	F_0_TO_7		:	STD_LOGIC;
SIGNAL	F_0_TO_7_STD:	STD_LOGIC_VECTOR (2  DOWNTO 0);

SIGNAL	F_8_TO_9		:	STD_LOGIC;
SIGNAL	F_10			:	STD_LOGIC;


SIGNAL	F_8_TO_11	:	STD_LOGIC;
SIGNAL	F_12_TO_13	:	STD_LOGIC;



SIGNAL	COUNTER_RAM			:	NATURAL RANGE      0   TO 327679 :=0;



SIGNAL	BUFGCLK200M	:	STD_LOGIC;

SIGNAL	CLK200M		:	STD_LOGIC;
SIGNAL	CLK100M		:	STD_LOGIC;
SIGNAL	CNT200M		:	STD_LOGIC_VECTOR (2  DOWNTO 0):="000";


SIGNAL	CLK_100_200M:	STD_LOGIC;
SIGNAL	CLK_100_200M_BUFG:	STD_LOGIC;

SIGNAL	CLK200M_NEW	:	STD_LOGIC;
SIGNAL	CLK200M_NEW_BUFG	:	STD_LOGIC;

SIGNAL	CLK400M	:	STD_LOGIC;
SIGNAL	CLK400M_BUFG	:	STD_LOGIC;


SIGNAL	CLK200M_END	:	STD_LOGIC;
--SIGNAL	CLK200M_END_BUFG	:	STD_LOGIC;


SIGNAL	CNT400M		:	STD_LOGIC_VECTOR (3  DOWNTO 0);



SIGNAL	BLCK_PRCH_H	:	STD_LOGIC;
SIGNAL	BLCK_PRCH_V	:	STD_LOGIC;






--SIGNAL	AVANCE		:	NATURAL RANGE 0 TO 1;
--SIGNAL	AVANCE_LINE	:	STD_LOGIC_VECTOR (18  DOWNTO 0):=(OTHERS=>'0');
--SIGNAL	AVANCE_PIXEL:	STD_LOGIC_VECTOR (9  DOWNTO 0):=(OTHERS=>'0');


TYPE SKDPARAMETER IS ARRAY (0 TO 2, 0 TO 1) OF STD_LOGIC_VECTOR (13 DOWNTO 0);
CONSTANT excellent: SKDPARAMETER:=( ("00100111100001","00010010111100"),
											   ("10011011000011","00010110101110"),
												("00111101010011","00010010001101") );


TYPE PIXEL IS ARRAY (0 TO 2) OF STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL PIXEL_DATA: PIXEL;

SIGNAL R_1000: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL G_1000: STD_LOGIC_VECTOR (21 DOWNTO 0);

SIGNAL G_MAXV1: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL G_MINV1: STD_LOGIC_VECTOR (21 DOWNTO 0);

SIGNAL B_MAXV2: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL B_MINV2: STD_LOGIC_VECTOR (21 DOWNTO 0);

SIGNAL B_MAXV3: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL B_MINV3: STD_LOGIC_VECTOR (21 DOWNTO 0);





SIGNAL	R_BIT_CMPL	:	STD_LOGIC;
SIGNAL	G_BIT_CMPL	:	STD_LOGIC;
SIGNAL	B_BIT_CMPL	:	STD_LOGIC;


SIGNAL	IS_SKIN		:	BOOLEAN;
SIGNAL	IS_SKIN_CONV:	BOOLEAN;
SIGNAL	SKINVECTOR	:	STD_LOGIC_VECTOR (7 DOWNTO 0);




SIGNAL	X			:	NATURAL RANGE      0   TO 1023:=0;
SIGNAL	Y			:	NATURAL RANGE      0   TO 511:=0;


--SIGNAL	LINE_CUR	:	NATURAL RANGE      0   TO 307200:=0;



SIGNAL	COLOR_MARK_BIT	:	STD_LOGIC;
SIGNAL	COLOR_MARK_BIT1:	STD_LOGIC;
SIGNAL	MARK_BIT_X		:	STD_LOGIC;
SIGNAL	MARK_BIT_Y		:	STD_LOGIC;

SIGNAL	COLOR_MARK		:	STD_LOGIC_VECTOR (7  DOWNTO 0);
SIGNAL	COLOR_MARK_NOT	:	STD_LOGIC_VECTOR (7  DOWNTO 0);




BEGIN
	RED	<=	(COLOR(7 DOWNTO 5) AND ZERO_COLOR(7 DOWNTO 5))	WHEN	NORM_NEGA	ELSE
				(NOT COLOR(7 DOWNTO 5) AND ZERO_COLOR(7 DOWNTO 5));
	
	GRN	<=	(COLOR(4 DOWNTO 2) AND ZERO_COLOR(4 DOWNTO 2))	WHEN	NORM_NEGA	ELSE
				(NOT COLOR(4 DOWNTO 2) AND ZERO_COLOR(4 DOWNTO 2));
	
	BLUE	<=	(COLOR(1 DOWNTO 0) AND ZERO_COLOR(1 DOWNTO 0))	WHEN	NORM_NEGA	ELSE
				(NOT COLOR(1 DOWNTO 0) AND ZERO_COLOR(1 DOWNTO 0));
	

	
	
	
	R_BIT_CMPL	<=	COLOR_RED(5) AND 
						COLOR_RED(4) AND 
						COLOR_RED(3) AND 
						COLOR_RED(2) AND 
						COLOR_RED(1) AND 
						COLOR_RED(0);
	PIXEL_DATA(0)	<=	COLOR_RED&(R_BIT_CMPL&R_BIT_CMPL);
	
	
	
	G_BIT_CMPL	<=	COLOR_GREEN(5) AND 
						COLOR_GREEN(4) AND 
						COLOR_GREEN(3) AND 
						COLOR_GREEN(2) AND 
						COLOR_GREEN(1) AND 
						COLOR_GREEN(0);
	PIXEL_DATA(1)	<=	COLOR_GREEN&(G_BIT_CMPL&G_BIT_CMPL);
	
	
	
	
	
	
	B_BIT_CMPL	<=	COLOR_BLUE(3) AND 
						COLOR_BLUE(2) AND 
						COLOR_BLUE(1) AND 
						COLOR_BLUE(0);
	PIXEL_DATA(2)	<=	COLOR_BLUE&(B_BIT_CMPL&B_BIT_CMPL&B_BIT_CMPL&B_BIT_CMPL);
	
	
	
	
	R_1000<="00001111101000"*(PIXEL_DATA(0));
	G_1000<="00001111101000"*(PIXEL_DATA(1));

	G_MAXV1<=excellent(0,0)*(PIXEL_DATA(1));
	G_MINV1<=excellent(0,1)*(PIXEL_DATA(1));

	B_MAXV2<=excellent(1,0)*(PIXEL_DATA(2));
	B_MINV2<=excellent(1,1)*(PIXEL_DATA(2));

	B_MAXV3<=excellent(2,0)*(PIXEL_DATA(2));
	B_MINV3<=excellent(2,1)*(PIXEL_DATA(2));
	
	
	
	IS_SKIN	<=	(  ((R_1000>G_MINV1) AND (R_1000<G_MAXV1)) AND ((R_1000>B_MINV2) AND (R_1000<B_MAXV2)) AND 
												((G_1000>B_MINV3) AND (G_1000<B_MAXV3)) );
	
	
	IS_SKIN_CONV	<=	IS_SKIN OR (NOT SKD);
	SKINVECTOR	<=	(OTHERS=>TO_BIT(IS_SKIN_CONV));
												

	
	PROCESS (CLK25M)																  --VGA
	BEGIN
		IF (CLK25M'EVENT AND CLK25M='0') THEN
			
			IF POS_X_S(9)='1' AND
				NOT(POS_X_S(9)='1' AND POS_X_S(8)='1' AND POS_X_S(7)='1' ) AND
				POS_Y_S(8)='1' AND POS_Y_S(7)='1' AND POS_Y_S(6)='1' THEN
				
				MARK_BIT_X	<=	'1';
				MARK_BIT_Y	<=	'1';
			ELSE
				MARK_BIT_X	<=	'0';
				MARK_BIT_Y	<=	'0';
			END IF;
			
			
		END IF;
	END PROCESS;
	
	COLOR_MARK_BIT1	<=	COLOR_MARK_BIT AND MARK_BIT_X AND MARK_BIT_Y;
	
	--MARK_BIT_X	<=	POS_X_S(9);
	--MARK_BIT_Y	<=	POS_Y_S(8) AND POS_Y_S(7) AND POS_Y_S(6);--"111000000";
		
	COLOR_MARK	<=	(OTHERS=>(COLOR_MARK_BIT1 AND TO_BIT(MARK)));
	COLOR_MARK_NOT	<=	(OTHERS=>(NOT TO_BIT(MARK) OR NOT(MARK_BIT_X AND MARK_BIT_Y)));
			
			
	COLOR_MARK_BIT	<=	BY_ADRIAN_C_MARK( CONV_INTEGER((POS_Y_S(4 DOWNTO 0))) )( CONV_INTEGER(POS_X_S(6 DOWNTO 0)) );
	
	
	COLOR	<=	((((COLOR_16_BITS OR COLOR_8_BITS) AND SKINVECTOR) XOR COLOR_LETTER) AND 
				COLOR_MARK_NOT) OR COLOR_MARK;-- AND ZERO_COLOR;
	
	
	
	
	CNT_RAM_POS	<=	COUNTER_RAM;

	VS <= NOT TO_BIT(	(COUNTER_V<2) );
	HS <= NOT TO_BIT(	(COUNTER_H<96) );
	
	
----------------------------------------------------------------------------------------------------------------------
	--HORIZONTAL.
	BLCK_PRCH_H	<=	TO_BIT( (COUNTER_H<144 OR COUNTER_H>783) );
--	BLCK_PRCH_H	<=	( (NOT COUNTER_H(9)) AND (NOT COUNTER_H(8)) AND
--						NOT( COUNTER_H(7) AND ( COUNTER_H(6) OR COUNTER_H(5) OR COUNTER_H(4) ) )   )	OR
--						( COUNTER_H(9) AND COUNTER_H(8) AND  COUNTER_H(4) );
	--VERTICAL.
	BLCK_PRCH_V	<=	TO_BIT( (COUNTER_V<31  OR COUNTER_V>510) );
--	BLCK_PRCH_V	<=	( COUNTER_V(9) OR ( COUNTER_V(8) AND COUNTER_V(7) AND COUNTER_V(6) AND	--510
--													COUNTER_V(5) AND COUNTER_V(4) AND COUNTER_V(3)	) )	OR
--						( ( (NOT COUNTER_V(9)) AND (NOT COUNTER_V(8)) AND (NOT COUNTER_V(7)) AND (NOT COUNTER_V(6)) AND
--							(NOT COUNTER_V(5))) AND 
--							( COUNTER_V(4) OR COUNTER_V(3) OR COUNTER_V(2) OR COUNTER_V(1) OR ( NOT COUNTER_V(0)) ) );
--	AREA_NEGRA <= ( (COUNTER_H<144) OR (COUNTER_H>783) OR 
--						 (COUNTER_V<31)  OR (COUNTER_V>510) );
	
	
	
	
	VGA_16_8_VECTOR<=	( OTHERS=>(NOT TO_BIT(VGA_16_8)) );
	
	COLOR_8_BITS	<=	(COLOR_RED(5 DOWNTO 3)&COLOR_GREEN(5 DOWNTO 3)&COLOR_BLUE(3 DOWNTO 2) ) AND VGA_16_8_VECTOR;
	COLOR_16_BITS	<=	(TOCOLORRED&TOCOLORGREEN&TOCOLORBLUE) AND (NOT VGA_16_8_VECTOR);
	
	
	ZERO_COLOR	<=	(OTHERS=> ( NOT (BLCK_PRCH_V OR BLCK_PRCH_H) ) );
	
	
	
	

	
	

	F_0_TO_7		<=	NOT CNT400M(3);
	F_0_TO_7_STD<=	(OTHERS=>F_0_TO_7);
	
	F_8_TO_9		<=	CNT400M(3) AND (NOT CNT400M(2)) AND (NOT CNT400M(1));
	
	F_10		<=	CNT400M(3) AND (NOT CNT400M(2))	AND CNT400M(1) AND ( NOT CNT400M(0) );
	
	TOCOLORRED	<=	( COLOR_RED(5 DOWNTO 3) 	 AND F_0_TO_7_STD )				OR
						( '0'&COLOR_RED(2 DOWNTO 1) AND '0'&F_8_TO_9&F_8_TO_9 )	OR
						( '0'&'0'&COLOR_RED(0) 		 AND '0'&'0'&F_10 );

	
	TOCOLORGREEN<=	( COLOR_GREEN(5 DOWNTO 3) 		AND F_0_TO_7_STD )			OR
						( '0'&COLOR_GREEN(2 DOWNTO 1) AND '0'&F_8_TO_9&F_8_TO_9 )OR
						( '0'&'0'&COLOR_GREEN(0) 		AND '0'&'0'&F_10 );

	
	
	F_8_TO_11	<=	CNT400M(3) AND (NOT CNT400M(2));
	F_12_TO_13	<=	CNT400M(3) AND CNT400M(2) AND (NOT CNT400M(1));
	
	TOCOLORBLUE	<=	(COLOR_BLUE(3 DOWNTO 2) AND F_0_TO_7_STD(1 DOWNTO 0) )	OR 
						( '0'&COLOR_BLUE(1) AND F_8_TO_11&F_8_TO_11)	OR
						( '0'&COLOR_BLUE(0) AND F_12_TO_13&F_12_TO_13);
	
	
	
	
	
	
	
	
	
-------------------------------------------------------------------------------------
	POS_X	<=	POS_X_S;
	POS_Y	<=	POS_Y_S;
	
	POS_X_S	<=	COUNTER_H-144;
	POS_Y_S	<=	COUNTER_V(8 DOWNTO 0)-31;
	
	X	<=	CONV_INTEGER(POS_X_S(9 DOWNTO ZOOM))*CONV_INTEGER( (NOT TO_BIT(COUNTER_H_CUR<145)));
	Y	<=	CONV_INTEGER(POS_Y_S(8 DOWNTO ZOOM));
	
	
	
	
	
	COUNTER_RAM	<=	( (X+MOVE_X) + 640*Y+640*MOVE_Y )*
						CONV_INTEGER( TO_BIT( (NOT(COUNTER_H_CUR>790 AND COUNTER_V_CUR>518)) ) );

-------------------------------------------------------------------------------------

	PROCESS (CLK25M)																  --VGA
	BEGIN
		IF (CLK25M'EVENT AND CLK25M='1') THEN
			COUNTER_H<=	COUNTER_H_CUR;
			COUNTER_V<=	COUNTER_V_CUR;
		END IF;
	END PROCESS;
	--
	PROCESS (COUNTER_H,COUNTER_V,COUNTER_H_CUR,COUNTER_V_CUR)
	BEGIN
		CASE	COUNTER_H	IS
			WHEN "11"&x"1F" =>
				COUNTER_H_CUR	<=	(OTHERS=>'0');
			WHEN OTHERS =>
				COUNTER_H_CUR	<=	COUNTER_H+1;
		END CASE;
		
		CASE	COUNTER_V	IS
			WHEN "10"&x"08" =>
				COUNTER_V_CUR	<=	(OTHERS=>'0');
			WHEN OTHERS =>
				IF COUNTER_H_CUR="00"&X"00" THEN
					COUNTER_V_CUR	<=	COUNTER_V+1;
				ELSE
					COUNTER_V_CUR	<=	COUNTER_V;
				END IF;
		END CASE;
	END PROCESS;
	
	
	
	
	
	
	
-------------------------------------------------------------------------------------
	DRIVERCLKDLL100:	clkDllCtrl PORT	MAP ( CLK50M , CLK100M  );
	DRIVERCLKDLL200:	clkDllCtrl PORT	MAP ( CLK100M , CLK200M );
	
   BUFG_INST1 : BUFG
   PORT MAP (
      O => BUFGCLK200M,   -- CLOCK BUFFER OUTPUT
      I => CLK200M -- CLOCK BUFFER INPUT
   );
	
-------------------------------------------------------------------------------------
	PROCESS (BUFGCLK200M)
	BEGIN
		IF (BUFGCLK200M'EVENT AND BUFGCLK200M='1') THEN
			CLK_100_200M	<=	NOT CLK_100_200M;
			CNT200M	<=	CNT200M+1;
		END IF;
	END PROCESS;
-------------------------------------------------------------------------------------
   BUFG_INST100_200 : BUFG
   PORT MAP (
      O => CLK_100_200M_BUFG,
      I => CLK_100_200M
   );
	
	
	
	DRIVERCLKDLL_100_200:	clkDllCtrl PORT MAP ( CLK_100_200M_BUFG , CLK200M_NEW );
   BUFG_INST200_NEW : BUFG
   PORT MAP (
      O => CLK200M_NEW_BUFG,
      I => CLK200M_NEW
   );
	
	
	
	
	DRIVERCLKDLL_200_NEW:	clkDllCtrl PORT MAP ( CLK200M_NEW_BUFG , CLK400M );
   BUFG_INST400 : BUFG
   PORT MAP (
      O => CLK400M_BUFG,
      I => CLK400M
   );
-------------------------------------------------------------------------------------
	PROCESS (CLK400M_BUFG)
	BEGIN
		IF (CLK400M_BUFG'EVENT AND CLK400M_BUFG='1') THEN
			CLK200M_END	<=	NOT CLK200M_END;
		END IF;
	END PROCESS;
	
	CLK25M	<=	NOT CNT200M(2);
	
	CNT400M	<=	CNT200M&(NOT CLK200M_END);
	
-------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------
--   BUFG_INST200_END : BUFG
--   PORT MAP (
--      O => CLK200M_END_BUFG,
--      I => CLK200M_END
--   );
--	PROCESS (CLK200M_END_BUFG)
--	BEGIN
--		IF (CLK200M_END_BUFG'EVENT AND CLK200M_END_BUFG='1') THEN
--			--CNT200M	<=	CNT200M+1;			
--		END IF;
--	END PROCESS;
	
--	PROCESS (CLK200M_END)
--	BEGIN
--		IF (CLK200M_END'EVENT AND CLK200M_END='1') THEN
--			CNT200M	<=	CNT200M+1;			
--		END IF;
--	END PROCESS;




END BEHAVIORAL;