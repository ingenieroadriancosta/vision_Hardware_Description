LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
-----------------------------------------------------
ENTITY BYTE2BCDALL IS
	PORT (   BYTE    		:	IN    STD_LOGIC_VECTOR (7  DOWNTO 0);
				DIGITO0   	:	OUT   NATURAL RANGE 0 TO 15;
				DIGITO1   	:	OUT   NATURAL RANGE 0 TO 15;
				DIGITO2   	:	OUT   NATURAL RANGE 0 TO 15
-----------------------------------------------------------------
         );
END BYTE2BCDALL;
-----------------------------------------------------
ARCHITECTURE BEHAVIORAL OF BYTE2BCDALL IS

SIGNAL	DU0			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU1			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU2			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU3			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU4			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU5			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );

SIGNAL	DD0			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD1			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD2			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );

SIGNAL	DC0			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );

BEGIN
	--UNIDADES.
	DU0	<=	'0'&BYTE(7 DOWNTO 5)	WHEN	(BYTE(7 DOWNTO 5)<5)	ELSE
				'0'&BYTE(7 DOWNTO 5)+3;
	DU1	<=	DU0(2 DOWNTO 0)&BYTE(4)	WHEN	( (DU0(2 DOWNTO 0)&BYTE(4))<5 )	ELSE
				DU0(2 DOWNTO 0)&BYTE(4)+3;
	DU2	<=	DU1(2 DOWNTO 0)&BYTE(3)	WHEN	( (DU1(2 DOWNTO 0)&BYTE(3))<5 )	ELSE
				DU1(2 DOWNTO 0)&BYTE(3)+3;
	DU3	<=	DU2(2 DOWNTO 0)&BYTE(2)	WHEN	( (DU2(2 DOWNTO 0)&BYTE(2))<5 )	ELSE
				DU2(2 DOWNTO 0)&BYTE(2)+3;
	DU4	<=	DU3(2 DOWNTO 0)&BYTE(1)	WHEN	( (DU3(2 DOWNTO 0)&BYTE(1))<5 )	ELSE
				DU3(2 DOWNTO 0)&BYTE(1)+3;
	DU5	<=	DU4(2 DOWNTO 0)&BYTE(0);
	
	--DECENAS.
	DD0	<=	'0'&DU0(3)&DU1(3)&DU2(3)	WHEN	( (DU0(3)&DU1(3)&DU2(3))<5 )	ELSE
				'0'&DU0(3)&DU1(3)&DU2(3)+3;
	DD1	<=	DD0(2)&DD0(1)&DD0(0)&DU3(3)	WHEN	( (DD0(2)&DD0(1)&DD0(0)&DU3(3))<5 )	ELSE
				DD0(2)&DD0(1)&DD0(0)&DU3(3)+3;
	DD2	<=	DD1(2)&DD1(1)&DD1(0)&DU4(3);
	
	--CENTENAS.
	DC0	<=	'0'&'0'&DD0(3)&DD1(3);
	
	
--	DIGITO0	<=	DU5;
--	DIGITO1	<=	DD2;
--	DIGITO2	<=	DC0;

	DIGITO0	<=	CONV_INTEGER(DU5);
	DIGITO1	<=	CONV_INTEGER(DD2);
	DIGITO2	<=	CONV_INTEGER(DC0);
END BEHAVIORAL;