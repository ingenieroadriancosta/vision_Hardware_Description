LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
-----------------------------------------------------
ENTITY WORD2BCD IS
	PORT (   VARWORD	:	IN    STD_LOGIC_VECTOR (15  DOWNTO 0);
				UNIDAD	:	OUT   STD_LOGIC_VECTOR (3  DOWNTO 0);
				DECENA	:	OUT   STD_LOGIC_VECTOR (3  DOWNTO 0);
				CENTENA	:	OUT   STD_LOGIC_VECTOR (3  DOWNTO 0)
-----------------------------------------------------------------
         );
END WORD2BCD;
-----------------------------------------------------
ARCHITECTURE BEHAVIORAL OF WORD2BCD IS

SIGNAL	DU0			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU1			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU2			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU3			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU4			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU5			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU6			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU7			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU8			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU9			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU10			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU11			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU12			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DU13			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );

SIGNAL	DD0			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD1			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD2			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD3			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD4			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD5			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD6			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD7			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD8			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD9			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
SIGNAL	DD10			:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );

SIGNAL	DC0			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
SIGNAL	DC1			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
SIGNAL	DC2			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
SIGNAL	DC3			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
SIGNAL	DC4			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
SIGNAL	DC5			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
SIGNAL	DC6			:	STD_LOGIC_VECTOR( 1 DOWNTO 0 );
SIGNAL	DC7			:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );



BEGIN
	--UNIDADES.
	DU0	<=	'0'&VARWORD(15 DOWNTO 13)	WHEN	(VARWORD(15 DOWNTO 13)<5)	ELSE
				'0'&VARWORD(15 DOWNTO 13)+3;
	DU1	<=	DU0(2 DOWNTO 0)&VARWORD(12)	WHEN	( (DU0(2 DOWNTO 0)&VARWORD(12))<5 )	ELSE
				DU0(2 DOWNTO 0)&VARWORD(12)+3;
	DU2	<=	DU1(2 DOWNTO 0)&VARWORD(11)	WHEN	( (DU1(2 DOWNTO 0)&VARWORD(11))<5 )	ELSE
				DU1(2 DOWNTO 0)&VARWORD(11)+3;
	DU3	<=	DU2(2 DOWNTO 0)&VARWORD(10)	WHEN	( (DU2(2 DOWNTO 0)&VARWORD(10))<5 )	ELSE
				DU2(2 DOWNTO 0)&VARWORD(10)+3;
	DU4	<=	DU3(2 DOWNTO 0)&VARWORD(9)	WHEN	( (DU3(2 DOWNTO 0)&VARWORD(9))<5 )	ELSE
				DU3(2 DOWNTO 0)&VARWORD(9)+3;
	DU5	<=	DU4(2 DOWNTO 0)&VARWORD(8)	WHEN	( (DU4(2 DOWNTO 0)&VARWORD(8))<5 )	ELSE
				DU4(2 DOWNTO 0)&VARWORD(8)+3;
	DU6	<=	DU5(2 DOWNTO 0)&VARWORD(7)	WHEN	( (DU5(2 DOWNTO 0)&VARWORD(7))<5 )	ELSE
				DU5(2 DOWNTO 0)&VARWORD(7)+3;
	DU7	<=	DU6(2 DOWNTO 0)&VARWORD(6)	WHEN	( (DU6(2 DOWNTO 0)&VARWORD(6))<5 )	ELSE
				DU6(2 DOWNTO 0)&VARWORD(6)+3;
	DU8	<=	DU7(2 DOWNTO 0)&VARWORD(5)	WHEN	( (DU7(2 DOWNTO 0)&VARWORD(5))<5 )	ELSE
				DU7(2 DOWNTO 0)&VARWORD(5)+3;
	DU9	<=	DU8(2 DOWNTO 0)&VARWORD(4)	WHEN	( (DU8(2 DOWNTO 0)&VARWORD(4))<5 )	ELSE
				DU8(2 DOWNTO 0)&VARWORD(4)+3;
	DU10	<=	DU9(2 DOWNTO 0)&VARWORD(3)	WHEN	( (DU9(2 DOWNTO 0)&VARWORD(3))<5 )	ELSE
				DU9(2 DOWNTO 0)&VARWORD(3)+3;
	DU11	<=	DU10(2 DOWNTO 0)&VARWORD(2)	WHEN	( (DU10(2 DOWNTO 0)&VARWORD(2))<5 )	ELSE
				DU10(2 DOWNTO 0)&VARWORD(2)+3;
	DU12	<=	DU11(2 DOWNTO 0)&VARWORD(1)	WHEN	( (DU11(2 DOWNTO 0)&VARWORD(1))<5 )	ELSE
				DU11(2 DOWNTO 0)&VARWORD(1)+3;
	DU13	<=	DU12(2 DOWNTO 0)&VARWORD(0);
	
	--DECENAS.
	DD0	<=	'0'&DU0(3)&DU1(3)&DU2(3)	WHEN	( (DU0(3)&DU1(3)&DU2(3))<5 )	ELSE
				'0'&DU0(3)&DU1(3)&DU2(3)+3;
	DD1	<=	DD0(2)&DD0(1)&DD0(0)&DU3(3)	WHEN	( (DD0(2)&DD0(1)&DD0(0)&DU3(3))<5 )	ELSE
				DD0(2)&DD0(1)&DD0(0)&DU3(3)+3;
	DD2	<=	DD1(2)&DD1(1)&DD1(0)&DU4(3)	WHEN	( (DD1(2)&DD1(1)&DD1(0)&DU4(3))<5 )	ELSE
				DD1(2)&DD1(1)&DD1(0)&DU4(3)+3;
	DD3	<=	DD2(2)&DD2(1)&DD2(0)&DU5(3)	WHEN	( (DD2(2)&DD2(1)&DD2(0)&DU5(3))<5 )	ELSE
				DD2(2)&DD2(1)&DD2(0)&DU5(3)+3;
	DD4	<=	DD3(2)&DD3(1)&DD3(0)&DU6(3)	WHEN	( (DD3(2)&DD3(1)&DD3(0)&DU6(3))<5 )	ELSE
				DD3(2)&DD3(1)&DD3(0)&DU6(3)+3;
	DD5	<=	DD4(2)&DD4(1)&DD4(0)&DU7(3)	WHEN	( (DD4(2)&DD4(1)&DD4(0)&DU7(3))<5 )	ELSE
				DD4(2)&DD4(1)&DD4(0)&DU7(3)+3;
	DD6	<=	DD5(2)&DD5(1)&DD5(0)&DU8(3)	WHEN	( (DD5(2)&DD5(1)&DD5(0)&DU8(3))<5 )	ELSE
				DD5(2)&DD5(1)&DD5(0)&DU8(3)+3;
	DD7	<=	DD6(2)&DD6(1)&DD6(0)&DU9(3)	WHEN	( (DD6(2)&DD6(1)&DD6(0)&DU9(3))<5 )	ELSE
				DD6(2)&DD6(1)&DD6(0)&DU9(3)+3;
	DD8	<=	DD7(2)&DD7(1)&DD7(0)&DU10(3)	WHEN	( (DD7(2)&DD7(1)&DD7(0)&DU10(3))<5 )	ELSE
				DD7(2)&DD7(1)&DD7(0)&DU10(3)+3;
	DD9	<=	DD8(2)&DD8(1)&DD8(0)&DU11(3)	WHEN	( (DD8(2)&DD8(1)&DD8(0)&DU11(3))<5 )	ELSE
				DD8(2)&DD8(1)&DD8(0)&DU11(3)+3;
	DD10	<=	DD9(2)&DD9(1)&DD9(0)&DU12(3);
	
	
	--CENTENAS.
	DC0	<=	DD0(3)&DD1(3)&DD2(3)	WHEN	( ('0'&DD0(3)&DD1(3)&DD2(3))<5 )	ELSE
				DD0(3)&DD1(3)&DD2(3)+3;
	DC1	<=	DC0(1)&DC0(0)&DD3(3)	WHEN	( (DC0(2)&DC0(1)&DC0(0)&DD3(3))<5 )	ELSE
				DC0(1)&DC0(0)&DD3(3)+3;
	DC2	<=	DC1(1)&DC1(0)&DD4(3)	WHEN	( (DC1(2)&DC1(1)&DC1(0)&DD4(3))<5 )	ELSE
				DC1(1)&DC1(0)&DD4(3)+3;
	DC3	<=	DC2(1)&DC2(0)&DD5(3)	WHEN	( (DC2(2)&DC2(1)&DC2(0)&DD5(3))<5 )	ELSE
				DC2(1)&DC2(0)&DD5(3)+3;
	DC4	<=	DC3(1)&DC3(0)&DD6(3)	WHEN	( (DC3(2)&DC3(1)&DC3(0)&DD6(3))<5 )	ELSE
				DC3(1)&DC3(0)&DD6(3)+3;
	DC5	<=	DC4(1)&DC4(0)&DD7(3)	WHEN	( (DC4(2)&DC4(1)&DC4(0)&DD7(3))<5 )	ELSE
				DC4(1)&DC4(0)&DD7(3)+3;
	DC6	<=	DC5(0)&DD8(3)	WHEN	( (DC5(2)&DC5(1)&DC5(0)&DD8(3))<5 )	ELSE
				DC5(0)&DD8(3)+3;
	DC7	<=	DC6(1)&DC6(0)&DD9(3);
	
	
	
	
	
	UNIDAD	<=	DU13;
	DECENA	<=	DD10;
	CENTENA	<=	'0'&DC7;
	

END BEHAVIORAL;