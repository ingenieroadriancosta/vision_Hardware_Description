LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--			|MAYOR_LEVELS|			|MINOR_LEVELS|
--       |            |       |            |
--R/G		|        2529|       |        1212|
--R/B		|        9923|       |        1454|
--B/G		|        3923|       |        1165|
PACKAGE MYPACKAGES IS
TYPE SKDPARAMETER IS ARRAY (0 TO 2, 0 TO 1) OF STD_LOGIC_VECTOR (13 DOWNTO 0);
CONSTANT EXCELLENT: SKDPARAMETER:=( ("00100111100001","00010010111100"),
											   ("10011011000011","00010110101110"),
												("00111101010011","00010010001101") );
TYPE PIXEL IS ARRAY (0 TO 2) OF STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL PIXEL_DATA_TX1: PIXEL;
SIGNAL PIXEL_DATA_RX1: PIXEL;

SIGNAL R_1000: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL G_1000: STD_LOGIC_VECTOR (21 DOWNTO 0);

SIGNAL G_MAXV1: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL G_MINV1: STD_LOGIC_VECTOR (21 DOWNTO 0);

SIGNAL B_MAXV2: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL B_MINV2: STD_LOGIC_VECTOR (21 DOWNTO 0);

SIGNAL B_MAXV3: STD_LOGIC_VECTOR (21 DOWNTO 0);
SIGNAL B_MINV3: STD_LOGIC_VECTOR (21 DOWNTO 0);

END MYPACKAGES;